VERSION 5.7 ;
NOWIREEXTENSIONATTERMINAL OFF ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

LAYER pwell
  TYPE NWELL ;
END pwell

LAYER nwell  
  TYPE NWELL ;
END nwell

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER li1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 12.8 ;
  CAPACITANCE CPERSQDIST 164.0 ;
  EDGECAPACITANCE 57.0 ;
END li1

LAYER mcon
  TYPE CUT ;
  SPACING 0.19 ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 52.4 ;
  EDGECAPACITANCE 28.7 ;
  
  MANUFACTURINGGRID 0.005 ;
  
  ANTENNADIFFAREA 400.0 ;
  ANTENNACUMROUTINGPLUSCUT ;
  ANTENNAGATEPLUSDIFF 350.0 ;
  ANTENNAAREAFACTOR 400.0 ;
END met1

LAYER via
  TYPE CUT ;
  SPACING 0.17 ;
  ENCLOSURE BELOW 0.055 0.085 ;
  ENCLOSURE ABOVE 0.055 0.085 ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 52.4 ;
  EDGECAPACITANCE 28.7 ;
  
  MANUFACTURINGGRID 0.005 ;
  
  ANTENNADIFFAREA 400.0 ;
  ANTENNACUMROUTINGPLUSCUT ;
  ANTENNAGATEPLUSDIFF 350.0 ;
  ANTENNAAREAFACTOR 400.0 ;
END met2

LAYER via2
  TYPE CUT ;
  SPACING 0.20 ;
  ENCLOSURE BELOW 0.065 0.065 ;
  ENCLOSURE ABOVE 0.065 0.065 ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.68 ;
  WIDTH 0.30 ;
  SPACING 0.30 ;
  RESISTANCE RPERSQ 0.047 ;
  CAPACITANCE CPERSQDIST 39.2 ;
  EDGECAPACITANCE 23.1 ;
  
  MANUFACTURINGGRID 0.005 ;
  
  ANTENNADIFFAREA 400.0 ;
  ANTENNACUMROUTINGPLUSCUT ;
  ANTENNAGATEPLUSDIFF 350.0 ;
  ANTENNAAREAFACTOR 400.0 ;
END met3

LAYER via3
  TYPE CUT ;
  SPACING 0.20 ;
  ENCLOSURE BELOW 0.065 0.065 ;
  ENCLOSURE ABOVE 0.065 0.065 ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.30 ;
  SPACING 0.30 ;
  RESISTANCE RPERSQ 0.047 ;
  CAPACITANCE CPERSQDIST 39.2 ;
  EDGECAPACITANCE 23.1 ;
  
  MANUFACTURINGGRID 0.005 ;
  
  ANTENNADIFFAREA 400.0 ;
  ANTENNACUMROUTINGPLUSCUT ;
  ANTENNAGATEPLUSDIFF 350.0 ;
  ANTENNAAREAFACTOR 400.0 ;
END met4

LAYER via4
  TYPE CUT ;
  SPACING 0.32 ;
  ENCLOSURE BELOW 0.19 0.19 ;
  ENCLOSURE ABOVE 0.19 0.19 ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.60 ;
  WIDTH 0.80 ;
  SPACING 0.80 ;
  RESISTANCE RPERSQ 0.029 ;
  CAPACITANCE CPERSQDIST 31.2 ;
  EDGECAPACITANCE 18.5 ;
  
  MANUFACTURINGGRID 0.005 ;
  
  ANTENNADIFFAREA 400.0 ;
  ANTENNACUMROUTINGPLUSCUT ;
  ANTENNAGATEPLUSDIFF 350.0 ;
  ANTENNAAREAFACTOR 400.0 ;
END met5

LAYER via5
  TYPE CUT ;
  SPACING 0.32 ;
  ENCLOSURE BELOW 0.19 0.19 ;
  ENCLOSURE ABOVE 0.19 0.19 ;
END via5

LAYER met6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.60 ;
  WIDTH 0.80 ;
  SPACING 0.80 ;
  RESISTANCE RPERSQ 0.029 ;
  CAPACITANCE CPERSQDIST 31.2 ;
  EDGECAPACITANCE 18.5 ;
  
  MANUFACTURINGGRID 0.005 ;
  
  ANTENNADIFFAREA 400.0 ;
  ANTENNACUMROUTINGPLUSCUT ;
  ANTENNAGATEPLUSDIFF 350.0 ;
  ANTENNAAREAFACTOR 400.0 ;
END met6

SITE unithd
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 2.72 ;
END unithd

SITE unithd_16t
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 2.72 ;
END unithd_16t

MACRO sakemono90_fd_sc_hd__nand2_1
  CLASS CORE ;
  FOREIGN sakemono90_fd_sc_hd__nand2_1 0.0 0.0 ;
  ORIGIN 0.0 0.0 ;
  SIZE 0.92 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 0.725 1.405 ;
    END
  END A
  
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.405 1.405 ;
    END
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.575 0.425 1.905 ;
    END
  END Y

  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.720 ;
    END
  END VPWR

  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.000 0.920 0.240 ;
    END
  END VGND

  OBS
    LAYER li1 ;
      RECT 0.00 0.24 0.92 1.07 ;
      RECT 0.00 1.41 0.92 2.48 ;
  END

END sakemono90_fd_sc_hd__nand2_1

MACRO sakemono90_fd_sc_hd__nor2_1
  CLASS CORE ;
  FOREIGN sakemono90_fd_sc_hd__nor2_1 0.0 0.0 ;
  ORIGIN 0.0 0.0 ;
  SIZE 0.92 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 0.725 1.405 ;
    END
  END A
  
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.405 1.405 ;
    END
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.575 0.425 1.905 ;
    END
  END Y

  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.720 ;
    END
  END VPWR

  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.000 0.920 0.240 ;
    END
  END VGND

  OBS
    LAYER li1 ;
      RECT 0.00 0.24 0.92 1.07 ;
      RECT 0.00 1.41 0.92 2.48 ;
  END

END sakemono90_fd_sc_hd__nor2_1

MACRO sakemono90_fd_sc_hd__and2_1
  CLASS CORE ;
  FOREIGN sakemono90_fd_sc_hd__and2_1 0.0 0.0 ;
  ORIGIN 0.0 0.0 ;
  SIZE 1.38 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 0.725 1.405 ;
    END
  END A
  
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.405 1.405 ;
    END
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.575 1.355 1.905 ;
    END
  END Y

  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.720 ;
    END
  END VPWR

  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.000 1.380 0.240 ;
    END
  END VGND

  OBS
    LAYER li1 ;
      RECT 0.00 0.24 1.38 1.07 ;
      RECT 0.00 1.41 0.73 2.48 ;
      RECT 1.05 1.41 1.38 2.48 ;
  END

END sakemono90_fd_sc_hd__and2_1

MACRO sakemono90_fd_sc_hd__or2_1
  CLASS CORE ;
  FOREIGN sakemono90_fd_sc_hd__or2_1 0.0 0.0 ;
  ORIGIN 0.0 0.0 ;
  SIZE 1.38 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 0.725 1.405 ;
    END
  END A
  
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.405 1.405 ;
    END
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.575 1.355 1.905 ;
    END
  END Y

  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.720 ;
    END
  END VPWR

  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.000 1.380 0.240 ;
    END
  END VGND

  OBS
    LAYER li1 ;
      RECT 0.00 0.24 1.38 1.07 ;
      RECT 0.00 1.41 0.73 2.48 ;
      RECT 1.05 1.41 1.38 2.48 ;
  END

END sakemono90_fd_sc_hd__or2_1

END LIBRARY