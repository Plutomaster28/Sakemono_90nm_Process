VERSION 5.7 ;
NOWIREEXTENSIONATTERMINAL OFF ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

LAYER pwell
  TYPE NWELL ;
END pwell

LAYER nwell  
  TYPE NWELL ;
END nwell

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER li1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 12.8 ;
  CAPACITANCE CPERSQDIST 164.0 ;
  EDGECAPACITANCE 57.0 ;
END li1

LAYER mcon
  TYPE CUT ;
  SPACING 0.19 ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 52.4 ;
  EDGECAPACITANCE 28.7 ;
  
  MANUFACTURINGGRID 0.005 ;
  
  ANTENNADIFFAREA 400.0 ;
  ANTENNACUMROUTINGPLUSCUT ;
  ANTENNAGATEPLUSDIFF 350.0 ;
  ANTENNAAREAFACTOR 400.0 ;
END met1

LAYER via
  TYPE CUT ;
  SPACING 0.17 ;
  ENCLOSURE BELOW 0.055 0.085 ;
  ENCLOSURE ABOVE 0.055 0.085 ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 52.4 ;
  EDGECAPACITANCE 28.7 ;
  
  MANUFACTURINGGRID 0.005 ;
  
  ANTENNADIFFAREA 400.0 ;
  ANTENNACUMROUTINGPLUSCUT ;
  ANTENNAGATEPLUSDIFF 350.0 ;
  ANTENNAAREAFACTOR 400.0 ;
END met2

SITE unithd
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 2.72 ;
END unithd

SITE unithd_16t
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 2.72 ;
END unithd_16t

MACRO sakemono90_fd_sc_hd__buf_1
  CLASS CORE ;
  FOREIGN sakemono90_fd_sc_hd__buf_1 0.0 0.0 ;
  ORIGIN 0.0 0.0 ;
  SIZE 1.38 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.405 1.405 ;
    END
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.575 1.355 1.905 ;
    END
  END X

  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.720 ;
    END
  END VPWR

  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.000 1.380 0.240 ;
    END
  END VGND

  OBS
    LAYER li1 ;
      RECT 0.00 0.24 1.38 1.07 ;
      RECT 0.00 1.41 0.60 2.48 ;
      RECT 0.85 1.41 1.38 2.48 ;
  END

END sakemono90_fd_sc_hd__buf_1

MACRO sakemono90_fd_sc_hd__buf_2
  CLASS CORE ;
  FOREIGN sakemono90_fd_sc_hd__buf_2 0.0 0.0 ;
  ORIGIN 0.0 0.0 ;
  SIZE 1.84 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.405 1.405 ;
    END
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.575 1.815 1.905 ;
    END
  END X

  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.720 ;
    END
  END VPWR

  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.000 1.840 0.240 ;
    END
  END VGND

  OBS
    LAYER li1 ;
      RECT 0.00 0.24 1.84 1.07 ;
      RECT 0.00 1.41 0.60 2.48 ;
      RECT 1.06 1.41 1.84 2.48 ;
  END

END sakemono90_fd_sc_hd__buf_2

MACRO sakemono90_fd_sc_hd__buf_4
  CLASS CORE ;
  FOREIGN sakemono90_fd_sc_hd__buf_4 0.0 0.0 ;
  ORIGIN 0.0 0.0 ;
  SIZE 2.30 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.405 1.405 ;
    END
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.575 2.275 1.905 ;
    END
  END X

  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.720 ;
    END
  END VPWR

  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.000 2.300 0.240 ;
    END
  END VGND

  OBS
    LAYER li1 ;
      RECT 0.00 0.24 2.30 1.07 ;
      RECT 0.00 1.41 0.60 2.48 ;
      RECT 1.52 1.41 2.30 2.48 ;
  END

END sakemono90_fd_sc_hd__buf_4

MACRO sakemono90_fd_sc_hd__buf_8
  CLASS CORE ;
  FOREIGN sakemono90_fd_sc_hd__buf_8 0.0 0.0 ;
  ORIGIN 0.0 0.0 ;
  SIZE 3.22 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.405 1.405 ;
    END
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.575 3.195 1.905 ;
    END
  END X

  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.720 ;
    END
  END VPWR

  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.000 3.220 0.240 ;
    END
  END VGND

  OBS
    LAYER li1 ;
      RECT 0.00 0.24 3.22 1.07 ;
      RECT 0.00 1.41 0.60 2.48 ;
      RECT 2.44 1.41 3.22 2.48 ;
  END

END sakemono90_fd_sc_hd__buf_8

MACRO sakemono90_fd_sc_hd__buf_16
  CLASS CORE ;
  FOREIGN sakemono90_fd_sc_hd__buf_16 0.0 0.0 ;
  ORIGIN 0.0 0.0 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.405 1.405 ;
    END
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.735 1.575 5.035 1.905 ;
    END
  END X

  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.720 ;
    END
  END VPWR

  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.000 5.060 0.240 ;
    END
  END VGND

  OBS
    LAYER li1 ;
      RECT 0.00 0.24 5.06 1.07 ;
      RECT 0.00 1.41 0.60 2.48 ;
      RECT 4.28 1.41 5.06 2.48 ;
  END

END sakemono90_fd_sc_hd__buf_16

END LIBRARY